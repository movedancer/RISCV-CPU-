`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/05/25 15:55:29
// Design Name: 
// Module Name: instr_memory
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module instr_memory(
    input clka,
    input ena,
    input [31:0]addra,
    output wire [31:0]douta
    );
    reg [31:0] rf[1023:0];
    initial begin
//        rf[0]=32'h00000213;
//        rf[1]=32'h00000413;
//        rf[2]=32'h00100493;
//        rf[3]=32'h00f00513;
//        rf[4]=32'h00249893;
//        rf[5]=32'h00151913;
//        rf[6]=32'h00200813;
//        rf[7]=32'h00a22023;
//        rf[8]=32'h00022003;
//        rf[9]=32'h00880a13;
//        rf[10]=32'h41048833;
//        rf[11]=32'h00a84733;
//        rf[12]=32'h00976733;
//        rf[13]=32'hfe000de3;
//        rf[14]=32'h00000000;
//        rf[15]=32'h00000000;
//���ָ��
//        rf[0]=32'h03106093;        
//        rf[1]=32'h00209093;        
//        rf[2]=32'h01506113;        
//        rf[3]=32'h00211113;        
//        rf[4]=32'h0220a1b3;   
//����ָ�����
//          rf[0]=32'h01006093;
//          rf[1]=32'h00209093;    
//          rf[2]=32'h0100e093;        
//          rf[3]=32'h01006113;        
//          rf[4]=32'h00211113;        
//          rf[5]=32'h00116113;        
//          rf[6]=32'h00006193;        
//          rf[7]=32'h001101b3;        
//          rf[8]=32'h00006193;        
//          rf[9]=32'h403081b3;        
//          rf[10]=32'h402181b3;        
//          rf[11]=32'h00218193;        
//          rf[12]=32'h00006193;       
//          rf[13]=32'h40018193;       
//          rf[14]=32'h00109093;       
//          rf[15]=32'h001101b3;       
//          rf[16]=32'h0ff06093;       
//          rf[17]=32'h01009093;       
//          rf[18]=32'h0000a133;       
//          rf[19]=32'h0000b133;       
//          rf[20]=32'h4000a113;       
//          rf[21]=32'h4000a113; 
//Logic����
//            rf[0]=32'h001010b7;
//            rf[1]=32'h1010e093;           
//            rf[2]=32'h1000e113;          
//            rf[3]=32'h0020e0b3;           
//            rf[4]=32'h0fe0f193;           
//            rf[5]=32'h0011f0b3;           
//            rf[6]=32'h3000c213;           
//            rf[7]=32'h001240b3; 
//��λ����
//              rf[0]=32'h00404137;
//              rf[1]=32'h40416113;
//              rf[2]=32'h00706393;
//              rf[3]=32'h00506293;
//              rf[4]=32'h00806413;
//              rf[5]=32'h00811113;
//              rf[6]=32'h00711133;
//              rf[7]=32'h00815113;
//              rf[8]=32'h00515133;
//              rf[9]=32'h01311113;
//              rf[10]=32'h41015113;
//              rf[11]=32'h40815133;
//S_Linst����
//                rf[0]=32'h0ff06193;
//                rf[1]=32'h003021a3;
//                rf[2]=32'h0081d193;
//                rf[3]=32'h00302123;
//                rf[4]=32'h0dd06193;      
//                rf[5]=32'h003020a3;        
//                rf[6]=32'h0081d193;        
//                rf[7]=32'h00302023;        
//                rf[8]=32'h00300083;        
//                rf[9]=32'h00204083;        
//                rf[10]=32'h00000013;        
//                rf[11]=32'h0bb06193;        
//                rf[12]=32'h00302223;        
//                rf[13]=32'h00405083;        
//                rf[14]=32'h00401083;        
//                rf[15]=32'h09906193;        
//                rf[16]=32'h00302323;        
//                rf[17]=32'h00601083;        
//                rf[18]=32'h00605083;       
//                rf[19]=32'h04506193;        
//                rf[20]=32'h01019193;        
//                rf[21]=32'h0671e193;        
//                rf[22]=32'h00302423;       
//                rf[23]=32'h00802083;
//��֧����bht
//                rf[0]=32'h00000293;        
//                rf[1]=32'h00000313;        
//                rf[2]=32'h00000393;        
//                rf[3]=32'h00a00e13;        
//                rf[4]=32'h00138393;        
//                rf[5]=32'h00530333;
//                rf[6]=32'h00128293;
//                rf[7]=32'hffc29ce3;
//                rf[8]=32'h00000293;
//                rf[9]=32'hffc396e3;
//                rf[10]=32'h00130313;
//��֧����btb
//                rf[0]=32'h00000293;        
//                rf[1]=32'h00000313;        
//                rf[2]=32'h06500393;        
//                rf[3]=32'h00530333;
//                rf[4]=32'h00128293;
//                rf[5]=32'hfe729ce3;
//                rf[6]=32'h00130313;
//�ۺϲ��Ծ���˷�
                rf[0]=32'h00404713;
                rf[1]=32'h00404693;
                rf[2]=32'h00e696b3;
                rf[3]=32'h00004633;
                rf[4]=32'h00e69533;
                rf[5]=32'h00a505b3;
                rf[6]=32'h000042b3;
                rf[7]=32'h00004333;
                rf[8]=32'h00004e33;
                rf[9]=32'h000043b3;
                rf[10]=32'h00e29eb3;
                rf[11]=32'h007e8eb3;
                rf[12]=32'h00ae8eb3;
                rf[13]=32'h000eae83;
                rf[14]=32'h00e39f33;
                rf[15]=32'h006f0f33;
                rf[16]=32'h00bf0f33;
                rf[17]=32'h000f2f03;
                rf[18]=32'h01eefeb3;
                rf[19]=32'h01de0e33;
                rf[20]=32'h00438393;
                rf[21]=32'hfcd3cae3;
                rf[22]=32'h00e29eb3;
                rf[23]=32'h006e8eb3;
                rf[24]=32'h00ce8eb3;
                rf[25]=32'h01cea023;
                rf[26]=32'h00430313;
                rf[27]=32'hfad34ae3;
                rf[28]=32'h00428293;
                rf[29]=32'hfad2c4e3;
                rf[30]=32'h0000006f;
//�ۺϲ�������
//                  rf[0]=32'h10004693;        
//                  rf[1]=32'h00001137;        
//                  rf[2]=32'h00004533;        
//                  rf[3]=32'h000045b3;        
//                  rf[4]=32'hfff68613;         
//                  rf[5]=32'h00261613;         
//                  rf[6]=32'h008000ef;         
//                  rf[7]=32'h0000006f;
//                  rf[8]=32'h0cc5da63;        
//                  rf[9]=32'h0005e333;        
//                  rf[10]=32'h000663b3;        
//                  rf[11]=32'h006502b3;       
//                  rf[12]=32'h0002a283;        
//                  rf[13]=32'h04735263;        
//                  rf[14]=32'h00750e33;        
//                  rf[15]=32'h000e2e03;        
//                  rf[16]=32'h005e4663;        
//                  rf[17]=32'hffc38393;        
//                  rf[18]=32'hfedff06f;        
//                  rf[19]=32'h00650eb3;
//                  rf[20]=32'h01cea023;
//                  rf[21]=32'h02735263; 
//                  rf[22]=32'h00650e33; 
//                  rf[23]=32'h000e2e03; 
//                  rf[24]=32'h01c2c663; 
//                  rf[25]=32'h00430313; 
//                  rf[26]=32'hfedff06f; 
//                  rf[27]=32'h00750eb3; 
//                  rf[28]=32'h01cea023; 
//                  rf[29]=32'hfc7340e3; 
//                  rf[30]=32'h00650eb3; 
//                  rf[31]=32'h005ea023; 
//                  rf[32]=32'hffc10113; 
//                  rf[33]=32'h00112023; 
//                  rf[34]=32'hffc10113; 
//                  rf[35]=32'h00b12023; 
//                  rf[36]=32'hffc10113; 
//                  rf[37]=32'h00c12023; 
//                  rf[38]=32'hffc10113; 
//                  rf[39]=32'h00612023; 
//                  rf[40]=32'hffc30613; 
//                  rf[41]=32'hf7dff0ef; 
//                  rf[42]=32'h00012303; 
//                  rf[43]=32'h00410113; 
//                  rf[44]=32'h00012603; 
//                  rf[45]=32'h00410113; 
//                  rf[46]=32'h00012583; 
//                  rf[47]=32'hffc10113; 
//                  rf[48]=32'h00c12023; 
//                  rf[49]=32'hffc10113; 
//                  rf[50]=32'h00612023; 
//                  rf[51]=32'h00430593; 
//                  rf[52]=32'hf51ff0ef; 
//                  rf[53]=32'h00012303; 
//                  rf[54]=32'h00410113; 
//                  rf[55]=32'h00012603; 
//                  rf[56]=32'h00410113; 
//                  rf[57]=32'h00012583; 
//                  rf[58]=32'h00410113; 
//                  rf[59]=32'h00012083; 
//                  rf[60]=32'h00410113; 
//                  rf[61]=32'h00008067;
    end
 //   wire [31:0]data;
//    always@(posedge clka)begin
//        if(ena)begin
//            data<=rf[addra];
//        end
//    end
//    always@(*)begin
//        if(ena)begin
//            assign data=rf[addra];
//        end
//    end
    assign douta=(ena)?rf[addra]:32'b0;
//    assign douta=data;
endmodule
